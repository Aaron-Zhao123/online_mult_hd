library verilog;
use verilog.vl_types.all;
entity testbench_mult_hd is
end testbench_mult_hd;
